// DE0_CV_QSYS_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module DE0_CV_QSYS_tb (
	);

	wire         de0_cv_qsys_inst_clk_bfm_clk_clk;                            // DE0_CV_QSYS_inst_clk_bfm:clk -> [DE0_CV_QSYS_inst:clk_clk, DE0_CV_QSYS_inst_reset_bfm:clk]
	wire         sdram_my_partner_clk_bfm_clk_clk;                            // sdram_my_partner_clk_bfm:clk -> sdram_my_partner:clk
	wire   [3:0] de0_cv_qsys_inst_key_external_connection_bfm_conduit_export; // DE0_CV_QSYS_inst_key_external_connection_bfm:sig_export -> DE0_CV_QSYS_inst:key_external_connection_export
	wire         de0_cv_qsys_inst_pll_locked_export;                          // DE0_CV_QSYS_inst:pll_locked_export -> DE0_CV_QSYS_inst_pll_locked_bfm:sig_export
	wire         de0_cv_qsys_inst_sdram_wire_cs_n;                            // DE0_CV_QSYS_inst:sdram_wire_cs_n -> sdram_my_partner:zs_cs_n
	wire   [1:0] de0_cv_qsys_inst_sdram_wire_dqm;                             // DE0_CV_QSYS_inst:sdram_wire_dqm -> sdram_my_partner:zs_dqm
	wire         de0_cv_qsys_inst_sdram_wire_cas_n;                           // DE0_CV_QSYS_inst:sdram_wire_cas_n -> sdram_my_partner:zs_cas_n
	wire         de0_cv_qsys_inst_sdram_wire_ras_n;                           // DE0_CV_QSYS_inst:sdram_wire_ras_n -> sdram_my_partner:zs_ras_n
	wire         de0_cv_qsys_inst_sdram_wire_we_n;                            // DE0_CV_QSYS_inst:sdram_wire_we_n -> sdram_my_partner:zs_we_n
	wire  [12:0] de0_cv_qsys_inst_sdram_wire_addr;                            // DE0_CV_QSYS_inst:sdram_wire_addr -> sdram_my_partner:zs_addr
	wire         de0_cv_qsys_inst_sdram_wire_cke;                             // DE0_CV_QSYS_inst:sdram_wire_cke -> sdram_my_partner:zs_cke
	wire  [15:0] de0_cv_qsys_inst_sdram_wire_dq;                              // [] -> [DE0_CV_QSYS_inst:sdram_wire_dq, sdram_my_partner:zs_dq]
	wire   [1:0] de0_cv_qsys_inst_sdram_wire_ba;                              // DE0_CV_QSYS_inst:sdram_wire_ba -> sdram_my_partner:zs_ba
	wire         de0_cv_qsys_inst_reset_bfm_reset_reset;                      // DE0_CV_QSYS_inst_reset_bfm:reset -> DE0_CV_QSYS_inst:reset_reset_n

	DE0_CV_QSYS de0_cv_qsys_inst (
		.clk_clk                        (de0_cv_qsys_inst_clk_bfm_clk_clk),                            //                     clk.clk
		.clk_sdram_clk                  (),                                                            //               clk_sdram.clk
		.key_external_connection_export (de0_cv_qsys_inst_key_external_connection_bfm_conduit_export), // key_external_connection.export
		.pll_locked_export              (de0_cv_qsys_inst_pll_locked_export),                          //              pll_locked.export
		.reset_reset_n                  (de0_cv_qsys_inst_reset_bfm_reset_reset),                      //                   reset.reset_n
		.sdram_wire_addr                (de0_cv_qsys_inst_sdram_wire_addr),                            //              sdram_wire.addr
		.sdram_wire_ba                  (de0_cv_qsys_inst_sdram_wire_ba),                              //                        .ba
		.sdram_wire_cas_n               (de0_cv_qsys_inst_sdram_wire_cas_n),                           //                        .cas_n
		.sdram_wire_cke                 (de0_cv_qsys_inst_sdram_wire_cke),                             //                        .cke
		.sdram_wire_cs_n                (de0_cv_qsys_inst_sdram_wire_cs_n),                            //                        .cs_n
		.sdram_wire_dq                  (de0_cv_qsys_inst_sdram_wire_dq),                              //                        .dq
		.sdram_wire_dqm                 (de0_cv_qsys_inst_sdram_wire_dqm),                             //                        .dqm
		.sdram_wire_ras_n               (de0_cv_qsys_inst_sdram_wire_ras_n),                           //                        .ras_n
		.sdram_wire_we_n                (de0_cv_qsys_inst_sdram_wire_we_n)                             //                        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) de0_cv_qsys_inst_clk_bfm (
		.clk (de0_cv_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm de0_cv_qsys_inst_key_external_connection_bfm (
		.sig_export (de0_cv_qsys_inst_key_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 de0_cv_qsys_inst_pll_locked_bfm (
		.sig_export (de0_cv_qsys_inst_pll_locked_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) de0_cv_qsys_inst_reset_bfm (
		.reset (de0_cv_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (de0_cv_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_sdram_partner_module sdram_my_partner (
		.clk      (sdram_my_partner_clk_bfm_clk_clk),  //     clk.clk
		.zs_dq    (de0_cv_qsys_inst_sdram_wire_dq),    // conduit.dq
		.zs_addr  (de0_cv_qsys_inst_sdram_wire_addr),  //        .addr
		.zs_ba    (de0_cv_qsys_inst_sdram_wire_ba),    //        .ba
		.zs_cas_n (de0_cv_qsys_inst_sdram_wire_cas_n), //        .cas_n
		.zs_cke   (de0_cv_qsys_inst_sdram_wire_cke),   //        .cke
		.zs_cs_n  (de0_cv_qsys_inst_sdram_wire_cs_n),  //        .cs_n
		.zs_dqm   (de0_cv_qsys_inst_sdram_wire_dqm),   //        .dqm
		.zs_ras_n (de0_cv_qsys_inst_sdram_wire_ras_n), //        .ras_n
		.zs_we_n  (de0_cv_qsys_inst_sdram_wire_we_n)   //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (143000000),
		.CLOCK_UNIT (1)
	) sdram_my_partner_clk_bfm (
		.clk (sdram_my_partner_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
